`include "uvm_macros.svh"
import uvm_pkg::*;

`include "tb/interface.sv"
`include "env/agent/transaction.sv"
`include "env/agent/sequencer.sv"
`include "env/agent/sequence.sv"
`include "env/agent/driver.sv"
`include "env/agent/monitor.sv"
`include "env/scoreboard.sv"
`include "env/env.sv"
`include "test/test.sv"

module top;
    bit clk;
    bit reset;
    
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // clock period 10ns
    end
    
    // Reset signal
    initial begin
        reset = 1;
        repeat(5) @(posedge clk);
        reset = 0;
    end
    
    // Interface instantiation
    if intf(.clk(clk), .reset(reset));
    
    // DUT instantiation
    RISCVPipelined dut(
        .clk(clk),
        .reset(reset)
    );
    
    // Todo: 
    //  1. What exactly signal are we trying to get from the DUT for monitor
    //  2. What exactly signal are we passing into the DUT (basically just clk and rst)
    assign intf.monitor_pc = dut.PC_F;
    assign intf.monitor_instr = dut.instruction_F;
    assign intf.monitor_result = dut.result_W;
    
    initial begin
        // Register interface with UVM config database
        uvm_config_db#(virtual if)::set(null, "*", "vif", intf);

        // Need to specify the running test name here 
        // or in the command line when simulation
        run_test();
    end
    
    // Dumping waveform (optional)
    // initial begin
    //     $dumpfile("dump.vcd");
    //     $dumpvars(0, top);
    // end
endmodule